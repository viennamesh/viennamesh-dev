--  GEOM PARTITION : partition algorithm
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : Partition_Inter2d.cdl
--  Author : Benedicte MARTIN
--  Module : GEOM

class Inter2d from Partition 

	---Purpose: Computes the intersections between edges on a face
	--          stores result is SD as AsDes from BRepAlgo.

uses
    AsDes               from BRepAlgo,
    Edge                from TopoDS,
    Face                from TopoDS,
    Vertex              from TopoDS,
    MapOfShape          from TopTools,
    Real                from Standard,
    ListOfShape         from TopTools

is
    CompletPart2d(myclass ; AsDes : mutable AsDes from BRepAlgo;
                            F     :         Face  from TopoDS;
                            NewEdges :      MapOfShape from TopTools);
		      
      	---Purpose: Computes the intersections between the edges stored
      	--          is AsDes as descendants of <F> . Intersections is computed
      	--          between two edges if one of them is bound in NewEdges.


    FindEndVertex(myclass; VertList : ListOfShape from TopTools;
                           f,l      : Real        from Standard;
                           E        : Edge        from TopoDS;
                           First    : out Boolean from Standard;
                           DU       : out Real    from Standard)
        returns Vertex from TopoDS;
    ---Purpose: Returns a vertex  from  <VertList> having parameter on
    --          <E> most close  to  <f>  or  <l>.  <First>  is True if
    --          found vertex is closer  to <f>. <DU> returns parameter
    --          difference.
    
    AddVonE(myclass; V : Vertex from TopoDS;
                     E1,E2 : Edge from TopoDS;
                     AsDes : mutable AsDes from BRepAlgo;
                     F: Face from TopoDS)
        returns Vertex from TopoDS;
        ---Purpose: Put V in AsDes as intersection of E1 and E2.
        --          Check that vertex equal to V already exists on one
        --          of edges, in  such  a  case,  V  is  not added but
        --          existing vertex is updated to  be on E1 and E2 and
        --          is returned insead of V.
        --          Optional F is a face  E1  and  E2  are on. If F is
        --          provided, it is used  to  find  new vertices on E1
        --          and E2 resulting from intersection of new edges on
        --          the two  other  faces  the  F  interferes with and
        --          through which E1 and  E2  pass  too. This helps to
        --          avoid small edges.


    GetTolerance(myclass; theV : Vertex from TopoDS;
                          theU : Real from Standard;
                          theE : Edge from TopoDS;
                          theAsDes : AsDes from BRepAlgo)
        returns Real from Standard;
        ---Purpose: Returns  tolerance  theV   must   have  atfer  its
        --          addition to theE with  theU parameter. theAsDes is
        --          used to find pcurves of theE

end Inter2d;

